module my_design();

endmodule:my_design
